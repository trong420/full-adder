*******************************************************************************
* CDL netlist
*
* Library : full_adder
* Top Cell Name: full_adder3
* View Name: schematic
* Netlist created: 20.May.2022 00:14:18
*******************************************************************************

*.SCALE METER
.GLOBAL vdd,vss

*******************************************************************************
* Library Name: full_adder
* Cell Name:    full_adder3
* View Name:    schematic
*******************************************************************************

*.SUBCKT full_adder3 B A Cin Cout S
*.PININFO Cout:O S:O B:I A:I Cin:I

M29 n17 n16 vss vss nch w=1.1u l=0.13u m=1
M24 n21 n6 vss vss nch w=1.1u l=0.13u m=1
M2 n13 A vss vss nch w=1.1u l=0.13u m=1
M20 n6 n1 vdd vdd pch w=1.1u l=0.13u m=1
M26 n17 n21 n19 vdd pch w=1.1u l=0.13u m=1
M27 Cout n17 vdd vdd pch w=1.1u l=0.13u m=1
M22 n5 n1 vss vss nch w=1.1u l=0.13u m=1
M14 n14 B vdd vdd pch w=1.1u l=0.13u m=1
M12 S n20 n1 vss nch w=1.1u l=0.13u m=1
M4 n1 B n13 vss nch w=1.1u l=0.13u m=1
M6 n1 n13 B vss nch w=1.1u l=0.13u m=1
M18 n16 n14 vss vss nch w=1.1u l=0.13u m=1
M17 n16 n14 vdd vdd pch w=1.1u l=0.13u m=1
M23 n21 n6 vdd vdd pch w=1.1u l=0.13u m=1
M28 n17 n21 vss vss nch w=1.1u l=0.13u m=1
M19 n6 Cin vdd vdd pch w=1.1u l=0.13u m=1
M9 S n1 Cin vdd pch w=1.1u l=0.13u m=1
M11 n1 Cin S vdd pch w=1.1u l=0.13u m=1
M16 n23 A vss vss nch w=1.1u l=0.13u m=1
M15 n14 B n23 vss nch w=1.1u l=0.13u m=1
M30 Cout n17 vss vss nch w=1.1u l=0.13u m=1
M25 n19 n16 vdd vdd pch w=1.1u l=0.13u m=1
M5 B A n1 vdd pch w=1.1u l=0.13u m=1
M21 n6 Cin n5 vss nch w=1.1u l=0.13u m=1
M3 n1 B A vdd pch w=1.1u l=0.13u m=1
M7 n20 Cin vdd vdd pch w=1.1u l=0.13u m=1
M8 n20 Cin vss vss nch w=1.1u l=0.13u m=1
M13 n14 A vdd vdd pch w=1.1u l=0.13u m=1
M1 n13 A vdd vdd pch w=1.1u l=0.13u m=1
M10 S n1 n20 vss nch w=1.1u l=0.13u m=1
*.ENDS

.END
