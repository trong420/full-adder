*******************************************************************************
* CDL netlist
*
* Library : full_adder
* Top Cell Name: full_adder3
* View Name: extracted
* Netlist created: 25.May.2022 17:35:25
*******************************************************************************

*.SCALE METER

*******************************************************************************
* Library Name: full_adder
* Cell Name:    full_adder3
* View Name:    extracted
*******************************************************************************

.SUBCKT full_adder3

M29 n6 n13 n0 n25 pch w=1.1e-06 l=1.3e-07 as=3.74e-13 ps=2.88e-06 ad=3.74e-13 pd=2.88e-06
M2 n9 n1 n12 n20 nch w=1.1e-06 l=1.3e-07 as=3.74e-13 ps=2.88e-06 ad=3.74e-13 pd=2.88e-06
M20 n14 n7 n9 n22 pch w=1.1e-06 l=1.3e-07 as=3.74e-13 ps=2.88e-06 ad=3.74e-13 pd=2.88e-06
M24 n0 n9 n10 n24 pch w=1.1e-06 l=1.3e-07 as=3.74e-13 ps=2.88e-06 ad=3.74e-13 pd=2.88e-06
M26 n0 n10 n16 n24 pch w=1.1e-06 l=1.3e-07 as=3.74e-13 ps=2.88e-06 ad=3.74e-13 pd=2.88e-06
M27 n0 n16 n13 n25 pch w=1.1e-06 l=1.3e-07 as=3.74e-13 ps=2.88e-06 ad=3.74e-13 pd=2.88e-06
M22 n18 n12 n2 n23 pch w=1.1e-06 l=1.3e-07 as=3.74e-13 ps=2.88e-06 ad=3.74e-13 pd=2.88e-06
M0 n5 n8 n1 n20 nch w=1.1e-06 l=1.3e-07 as=3.74e-13 ps=2.88e-06 ad=3.74e-13 pd=2.88e-06
M14 n6 n13 n5 n20 nch w=1.1e-06 l=1.3e-07 as=3.74e-13 ps=2.88e-06 ad=3.74e-13 pd=2.88e-06
M12 n13 n16 n5 n20 nch w=1.1e-06 l=1.3e-07 as=3.74e-13 ps=2.88e-06 ad=3.74e-13 pd=2.88e-06
M4 n9 n9 n14 n20 nch w=1.1e-06 l=1.3e-07 as=3.74e-13 ps=2.88e-06 ad=3.74e-13 pd=2.88e-06
M18 n0 n7 n9 n22 pch w=1.1e-06 l=1.3e-07 as=3.74e-13 ps=2.88e-06 ad=3.74e-13 pd=2.88e-06
M6 n5 n8 n3 n20 nch w=1.1e-06 l=1.3e-07 as=3.74e-13 ps=2.88e-06 ad=3.74e-13 pd=2.88e-06
M17 n9 n8 n12 n21 pch w=1.1e-06 l=1.3e-07 as=3.74e-13 ps=2.88e-06 ad=3.74e-13 pd=2.88e-06
M23 n0 n2 n4 n23 pch w=1.1e-06 l=1.3e-07 as=3.74e-13 ps=2.88e-06 ad=3.74e-13 pd=2.88e-06
M28 n13 n4 n17 n25 pch w=1.1e-06 l=1.3e-07 as=3.74e-13 ps=2.88e-06 ad=3.74e-13 pd=2.88e-06
M19 n7 n9 n14 n22 pch w=1.1e-06 l=1.3e-07 as=3.74e-13 ps=2.88e-06 ad=3.74e-13 pd=2.88e-06
M11 n16 n10 n5 n20 nch w=1.1e-06 l=1.3e-07 as=3.74e-13 ps=2.88e-06 ad=3.74e-13 pd=2.88e-06
M16 n8 n12 n9 n21 pch w=1.1e-06 l=1.3e-07 as=3.74e-13 ps=2.88e-06 ad=3.74e-13 pd=2.88e-06
M9 n5 n9 n15 n20 nch w=1.1e-06 l=1.3e-07 as=3.74e-13 ps=2.88e-06 ad=3.74e-13 pd=2.88e-06
M15 n0 n8 n1 n21 pch w=1.1e-06 l=1.3e-07 as=3.74e-13 ps=2.88e-06 ad=3.74e-13 pd=2.88e-06
M25 n19 n7 n10 n24 pch w=1.1e-06 l=1.3e-07 as=3.74e-13 ps=2.88e-06 ad=3.74e-13 pd=2.88e-06
M5 n14 n9 n9 n20 nch w=1.1e-06 l=1.3e-07 as=3.74e-13 ps=2.88e-06 ad=3.74e-13 pd=2.88e-06
M3 n5 n7 n9 n20 nch w=1.1e-06 l=1.3e-07 as=3.74e-13 ps=2.88e-06 ad=3.74e-13 pd=2.88e-06
M21 n0 n8 n2 n23 pch w=1.1e-06 l=1.3e-07 as=3.74e-13 ps=2.88e-06 ad=3.74e-13 pd=2.88e-06
M8 n5 n2 n4 n20 nch w=1.1e-06 l=1.3e-07 as=3.74e-13 ps=2.88e-06 ad=3.74e-13 pd=2.88e-06
M7 n3 n12 n2 n20 nch w=1.1e-06 l=1.3e-07 as=3.74e-13 ps=2.88e-06 ad=3.74e-13 pd=2.88e-06
M13 n13 n4 n11 n20 nch w=1.1e-06 l=1.3e-07 as=3.74e-13 ps=2.88e-06 ad=3.74e-13 pd=2.88e-06
M1 n1 n12 n9 n20 nch w=1.1e-06 l=1.3e-07 as=3.74e-13 ps=2.88e-06 ad=3.74e-13 pd=2.88e-06
M10 n10 n7 n15 n20 nch w=1.1e-06 l=1.3e-07 as=3.74e-13 ps=2.88e-06 ad=3.74e-13 pd=2.88e-06
.ENDS
